library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

-- substitua entity_template pela sua entidade

entity entity_template is 
  port();
end;

architecture arq of entity_template is

-- declare componentes e signals aqui

begin

  -- defina o comportamento aqui
end arq;
