LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;

ENTITY rom IS
  PORT (
    clk : IN STD_LOGIC;
    address : IN unsigned(6 DOWNTO 0);
    data : OUT unsigned(15 DOWNTO 0)
  );
END ENTITY;

ARCHITECTURE a_rom OF rom IS
  TYPE mem IS ARRAY (0 TO 127) OF unsigned(15 DOWNTO 0);
  CONSTANT content : mem := (

    ------------TESTE 19XXX (SELECIONA)------------
    0 => B"000000000_001_1001", --LU R1, 0x0000
    1 => B"010001011_000_1110", --LD A, 0x008B
    2 => B"000000000_001_0100", --ADD A, R1
    3 => B"000000000_001_0010", --MOV R1, A

    4 => B"000001100_010_1111", --LD R2, 0x000C  

    ------------TESTE 32 (SELECIONA)------------
    --0 => B"000000000_001_1001", --LU R1, 0x0000
    --1 => B"000100000_000_1110", --LD A, 0x0020
    --2 => B"000000000_001_0100", --ADD A, R1
    --3 => B"000000000_001_0010", --MOV R1, A

    --4 => B"000000110_010_1111", --LD R2, 0x0006    

    --Inicializa vetor com valores padroes
    5 => B"000000000_011_1111", --LD R3, 0
    6 => B"000000011_000_0111", --SW R0, R3
    7 => B"000000001_011_1111", --LD R3, 1
    8 => B"000000011_000_0111", --SW R0, R3

    9 => B"000000001_101_1111", --LD R5, 1
    10 => B"000000001_011_1111", --LD R3, 1
    11 => B"000000001_000_1110", --LD A, 1      : X
    12 => B"000000000_011_0100", --ADD A, R3
    13 => B"000000000_011_0010", --MOV R3, A
    14 => B"000000011_101_0111", --SW R5, R3
    15 => B"000000000_000_1101", --CLR Z
    16 => B"000000000_001_0011", --MOV A, R1
    17 => B"000000000_011_0101", --SUB A, R3
    18 => B"111111001_111_1100", --JB 7, X  / BNE X

    19 => B"011111111_111_1111", --LD R7, 0x00FF    <------ FLAG COMPLETED

    --Crivo algoritimo
    20 => B"000000001_011_1111", --LD R3, 1
    21 => B"000000001_000_1110", --LD A, 1                                   : Y
    22 => B"000000000_011_0100", --ADD A, R3
    23 => B"000000000_011_0010", --MOV R3, A
    24 => B"000000000_000_1101", --CLR Z
    25 => B"000000000_010_0011", --MOV A, R2
    26 => B"000000000_011_0101", --SUB A, R3
    27 => B"000010111_010_1100", --JB 2, END  /  BGT END
    28 => B"000000011_110_1000", --LW R6, R3
    29 => B"000000000_000_1101", --CLR Z
    30 => B"000000000_000_0011", --MOV A, R0
    31 => B"000000000_110_0101", --SUB A, R6
    32 => B"111110101_000_1100", --JB 0, Y  / BEQ Y
    33 => B"000000000_011_0011", --MOV A, R3
    34 => B"000000000_100_0010", --MOV R4, A
    35 => B"000000000_011_0011", --MOV A, R3                                  : Z
    36 => B"000000000_100_0100", --ADD A, R4
    37 => B"000000000_100_0010", --MOV R4, A
    38 => B"000000000_000_1101", --CLR Z
    39 => B"000000000_001_0011", --MOV A, R1
    40 => B"000000000_100_0101", --SUB R4, A
    41 => B"111101100_010_1100", --JB 2, Y  /  BGT Y
    42 => B"000000100_000_0111", --SW R0, R4
    43 => B"000100011_000_0001", --JMP Z

    50 => B"000000000_000_0000", --NOP                                        : END
    51 => B"011101101_111_1111", --LD R7, 0x00ED

    --Loop vetor crivo
    52 => B"000000000_011_1111", --LD R3, 0
    53 => B"000000001_000_1110", --LD A, 1                                    : loop
    54 => B"000000000_011_0100", --ADD A, R3
    55 => B"000000000_011_0010", --MOV R3, A
    56 => B"000000011_110_1000", --LW R6, R3
    57 => B"000000000_000_1101", --CLR Z
    58 => B"000000000_001_0011", --MOV A, R1
    59 => B"000000000_011_0101", --SUB A, R3
    60 => B"111111001_111_1100", --JB 7, loop  /  BNE loop

    --61 => B"001011101_000_0001", --JMP END2           <---- JUST IF 32

    --Loop verifica primo
    62 => B"001001010_001_1001", --LU R1, 0x004A                  <---- Primo a se verificar
    63 => B"011010000_000_1110", --LD A, 0x00D0
    --62 => B"001000101_001_1001", --LU R1, 0x0045                    <---- Primo a se verificar
    --63 => B"001111111_000_1110", --LD A, 0x007F

    64 => B"000000000_001_0100", --ADD A, R1
    65 => B"000000000_001_0010", --MOV R1, A

    66 => B"010001011_010_1111", --LD R2, 0x008B 

    67 => B"000000001_111_1111", --LD R7, 0x0001

    68 => B"000000001_011_1111", --LD R3, 1
    69 => B"000000001_000_1110", --LD A, 1                                   : Y2
    70 => B"000000000_011_0100", --ADD A, R3
    71 => B"000000000_011_0010", --MOV R3, A
    72 => B"000000000_000_1101", --CLR Z
    73 => B"000000000_010_0011", --MOV A, R2
    74 => B"000000000_011_0101", --SUB A, R3
    75 => B"000010010_010_1100", --JB 2, END2  /  BGT END2
    76 => B"000000011_110_1000", --LW R6, R3
    77 => B"000000000_000_1101", --CLR Z
    78 => B"000000000_000_0011", --MOV A, R0
    79 => B"000000000_110_0101", --SUB A, R6
    80 => B"111110101_000_1100", --JB 0, Y2  / BEQ Y2
    81 => B"000000000_011_0011", --MOV A, R3
    82 => B"000000000_100_0010", --MOV R4, A
    83 => B"000000000_011_0011", --MOV A, R3                                  : Z2
    84 => B"000000000_100_0100", --ADD A, R4
    85 => B"000000000_100_0010", --MOV R4, A
    86 => B"000000000_000_1101", --CLR Z
    87 => B"000000000_001_0011", --MOV A, R1
    88 => B"000000000_100_0101", --SUB R4, A
    89 => B"111101100_010_1100", --JB 2, Y2  /  BGT Y2
    90 => B"000000010_000_1100", --JB 0, NUMERO  /  BEQ NUMERO
    91 => B"001010011_000_0001", --JMP Z2

    92 => B"000000000_111_1111", --LD R7 0x0000                           :NUMERO
    93 => B"000000000_000_0000", --NOP                                      :END2
    OTHERS => (OTHERS => '0')
  );

  SIGNAL rom_data : unsigned(15 DOWNTO 0) := "0000000000000000";

BEGIN
  PROCESS (clk)
  BEGIN
    IF (rising_edge(clk)) THEN
      rom_data <= content(to_integer(address));
    END IF;
  END PROCESS;

  data <= rom_data;
END ARCHITECTURE;